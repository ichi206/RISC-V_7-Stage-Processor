package enums;

typedef enum {BYTE, HALFWORD, WORD} loadtype;

endpackage
